//design code
module add(
input [3:0] a,b,
output [4:0] y);
assign y=a+b;    
endmodule
