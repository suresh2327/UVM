//design code
module add(
input [3:0] a,b,
output [4:0] y);
assign y = a + b;    
<<<<<<< HEAD
endmodule
=======
endmodule
>>>>>>> f73e1af3ce620a02963dab30fe0aebe2bfa5eab0
